module DATAPATH(CLK,INST,REGDST,ALUSRC,ALUCONTROL,MEMWRITE,MEMREAD,MEMTOREG,OUT,REGWRITE);

input [25:0] INST;
output [31:0] OUT;
input CLK;
input REGDST,ALUSRC,MEMWRITE,MEMREAD,MEMTOREG,REGWRITE;
input [2:0] ALUCONTROL;
wire [31:0] RD1,RD2,ALURESULT,O_SIGNEXTEND,READDATA,WD;
wire [4:0] WR;

MUX_32_bit #(.WIDTH(5)) mux1(.OP(REGDST),.A(INST[20:16]),.B(INST[15:11]),.O(WR));

REGFILE REG1(.RWE(REGWRITE),.WA(WR),.WD(WD),.RA1(INST[25:21]),.RA2(INST[20:16]),.CLK(CLK),.RD1(RD1),.RD2(RD2));

wire [31:0] OM2;
MUX_32_bit #(.WIDTH(32)) mux2(.OP(ALUSRC),.A(RD2),.B(O_SIGNEXTEND),.O(OM2));

ALU ALU1(.A(RD1),.B(OM2),.O(ALURESULT),.OP(ALUCONTROL),.OF());

SRAM SRAM1(.CLK(CLK),.WE(MEMWRITE),.RE(MEMREAD),.WD(RD2),.RA(READDATA),.ADDRESS(ALURESULT));

SIGN_EXTEND SignEXTEND(.I(INST[15:0]),.O(O_SIGNEXTEND));

MUX_32_bit #(.WIDTH(32)) mux3(.OP(MEMTOREG),.A(ALURESULT),.B(READDATA),.O(WD));

assign OUT=WD;	
endmodule
