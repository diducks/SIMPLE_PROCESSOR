module Control_Unit(OP,REGDST,MEMREAD,MEMWRITE,MEMTOREG,ALUOP,ALUSRC,REGWRITE);

input [5:0] OP;
output reg REGDST,MEMREAD,MEMWRITE,MEMTOREG,ALUSRC,REGWRITE;
output reg [1:0] ALUOP;

always @(*)
		case(OP)
		1://add 
		begin
			ALUOP=2'd2;
			ALUSRC=1'b0;
			REGDST=1'b1;
			REGWRITE=1'b1;
			MEMREAD=1'b0;
			MEMWRITE=1'b0;
			MEMTOREG=1'b0;
		end
		3://sub
		begin
			ALUOP=2'd3;
			ALUSRC=1'b0;
			REGDST=1'b1;
			REGWRITE=1'b1;
			MEMREAD=1'b0;
			MEMWRITE=1'b0;
			MEMTOREG=1'b0;
		end
		5://and
		begin
			ALUOP=2'd0;
			ALUSRC=1'b0;
			REGDST=1'b1;
			REGWRITE=1'b1;
			MEMREAD=1'b0;
			MEMWRITE=1'b0;
			MEMTOREG=1'b0;
		end
		7://or
		begin
			ALUOP=2'd1;
			ALUSRC=1'b0;
			REGDST=1'b1;
			REGWRITE=1'b1;
			MEMREAD=1'b0;
			MEMWRITE=1'b0;
			MEMTOREG=1'b0;
		end
		4://lw
		begin
			ALUOP=2'd2;
			ALUSRC=1'b1;
			REGDST=1'b0;
			REGWRITE=1'b1;
			MEMREAD=1'b1;
			MEMWRITE=1'b0;
			MEMTOREG=1'b1;
		end
		2://sw
		begin
			ALUOP=2'd2;
			ALUSRC=1'b1;
			REGDST=1'b0;
			REGWRITE=1'b1;
			MEMREAD=1'b0;
			MEMWRITE=1'b1;
			MEMTOREG=1'b0;
		end
		default:
		begin
			ALUOP=2'dx;
			ALUSRC=1'bx;
			REGDST=1'bx;
			REGWRITE=1'bx;
			MEMREAD=1'bx;
			MEMWRITE=1'bx;
			MEMTOREG=1'bx;
		end
	endcase
endmodule