`timescale 1ns/100ps
module tb;
reg [31:0]INST;
reg CLK;
wire [31:0] OUT;
LAB07 uut(.INST(INST),.CLK(CLK),.OUT(OUT));
initial begin
#0 CLK=0;
end
initial begin
#0 INST=32'b000001_00010_00001_00001_00000000000;//add $1,$2,$1 
#1 $display("OUTPUT :%d",OUT);
#9 INST=32'b000001_00010_00011_00001_00000000000;//add $1,$2,$3
#10 INST=32'b000001_00100_00011_00010_00000000000;//add $2,$4,$3
#10 INST=32'b000011_00010_00011_00001_00000000000;//sub $1,$2,$3
#10 INST=32'b000100_00010_00011_0000000000000000;//lw $3,0($2);
#10 INST=32'b000010_00001_00010_0000000000000000;//sw $2,0($2);
#10 INST=32'b000111_00001_00010_0000000000000000;//or $2,0($2);
#10 INST=32'b000101_00001_00010_0000000000000000;//and $2,0($2);
end
always #5 begin 
#0 CLK=~CLK;
end
always #10 begin
#0 $display("OUTPUT :%d",OUT);
end
endmodule
