//module MUX_32_bit(OP,A,B,O);
//parameter WIDTH = 32;
//input [WIDTH-1:0] A,B;
//input OP;
//output reg [WIDTH-1:0] O;
//always @(*) begin
//O=(OP==0)?A:B;
//end
//endmodule
