module LAB07(INST,CLK,OUT);//,REGDST,ALUSRC,MEMWRITE,MEMREAD,MEMTOREG,REGWRITE);

input [31:0] INST;
input CLK;
output [31:0] OUT;

 wire REGDST,ALUSRC,MEMWRITE,MEMREAD,MEMTOREG,REGWRITE;
 wire [1:0] ALUOP;
 wire [2:0] ALUCONTROL;


DATAPATH DATAPATH1(.CLK(CLK),.INST(INST[25:0]),.REGDST(REGDST),.ALUSRC(ALUSRC),.ALUCONTROL(ALUCONTROL),.MEMWRITE(MEMWRITE),.MEMREAD(MEMREAD),.MEMTOREG(MEMTOREG),.OUT(OUT),.REGWRITE(REGWRITE));

Control_Unit Control_Unit1(.OP(INST[31:26]),.REGDST(REGDST),.MEMREAD(MEMREAD),.MEMWRITE(MEMWRITE),.MEMTOREG(MEMTOREG),.ALUOP(ALUOP),.ALUSRC(ALUSRC),.REGWRITE(REGWRITE));
Alu_control Alu_control1(.ALUOP(ALUOP),.ALUcontrol(ALUCONTROL));


endmodule
//000001_00000_00001_00010_00000000000 add $2,$1,$0
// thanh ghi $2 = 2 
//000001_00000_00010_00011_00000000000 add $3,$1,$2

